module CPU();

endmodule
